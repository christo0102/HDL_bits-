module top_module (
    input clk,
    input reset,
    input [7:0] d,
    output [7:0] q
);
    always @(negedge clk)begin
        if(reset)
            q<=6'd52;
        else
            q[7:0]<=d[7:0];
    end
endmodule
