module top_module ( input a, input b, output out );
    mod_a uut (a,b,out);
endmodule
